module parallel_txrx(
    output clock,
    input chip_select,
    inout [7:0] data
);

endmodule