`ifndef _parameters_vh_
`define _parameters_vh_
`define BAUD_RATE 460800
`define CLK_FREQUENCY 50000000
`endif